FUCK<1050>Arthur Dent<42>