1035604112