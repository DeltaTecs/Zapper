1.0;true;true;true;true;false