1.1;true;true;false;true;false