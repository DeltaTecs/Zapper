<24576>Arthur Dent<42>