Arthur Dent<42>fuck<0>jackpott<0>