Arthur Dent<42>