1.0;true;true;false;true;true;false;false