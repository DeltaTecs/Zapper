1.2;true;true;true;true;false