1.3;true;true;false;true;true