Arthur Dent<42