Da_BOSS<57856456>asd<57856456>name<57856456>Arthur Dent<42>Nigga<0>Nigga<0>Nigga<0>NIGGA<0>NIGA<0>