1035580583