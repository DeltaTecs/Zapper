1.0f;true;true;false;true;true;false;true