1035628308