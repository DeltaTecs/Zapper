1035628078