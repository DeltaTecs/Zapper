1.2;true;true;false;true;false