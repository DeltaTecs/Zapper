1035628170