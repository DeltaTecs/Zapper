1.0;true;true;false;true;false