1.25;true;true;false;true;false