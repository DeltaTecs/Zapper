Arthur Dent<42>DeezNutz<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>fuuuuuuuu<0>Name<0>awwwwwwwwwwwwwdwasdwa<0>wdasdawdasd<0>