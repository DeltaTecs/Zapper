1.0;true;true;false;false;false