trueBOIfalseBOIfalseBOItrueBOIfalseBOItrueBOIfalseBOIfalseBOIfalseBOIfalseBOItrue