1035628239