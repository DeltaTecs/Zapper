1035628331